module data_memory_tb();
	reg clk;
	reg we;
	reg a;

endmodule
